module UnicornPower (iGrayMem1,
							iGrayMem2
							);
							
input iGrayMem1;
input iGrayMem2;

							
endmodule